module m_and16 (
  input i_16bit_a,
  input i_16bit_b,
  output o_16bit_out
  )
