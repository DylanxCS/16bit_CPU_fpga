module m_not(
  input i_a,
  output o_out)
  
assign o_out = ~i_a;

endmodule
