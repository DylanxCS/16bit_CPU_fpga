module m_or (
  input i_a,
  input i_b,
  output o_out);

assign o_out = (i_a || i_b);
  
endmodule
