module m_not16 (
  input [15:0] i_16bit,
  output [15:0] o_16bit
  );
 
m_not bit1 (
 .i_a(i_16bit[0]),
 .o_out(o_16bit[0])
 );
 
m_not bit2 (
 .i_a(i_16bit[1]),
 .o_out(o_16bit[1])
 );
 
m_not bit3 (
 .i_a(i_16bit[2]),
 .o_out(o_16bit[2])
 );
 
m_not bit4 (
 .i_a(i_16bit[3]),
 .o_out(o_16bit[3])
 );
 
m_not bit5 (
 .i_a(i_16bit[4]),
 .o_out(o_16bit[4])
 );
 
m_not bit6 (
 .i_a(i_16bit[5]),
 .o_out(o_16bit[5])
 );
 
m_not bit7 (
 .i_a(i_16bit[6]),
 .o_out(o_16bit[6])
 );
 
m_not bit8 (
 .i_a(i_16bit[7]),
 .o_out(o_16bit[7])
 );
 
m_not bit9 (
 .i_a(i_16bit[8]),
 .o_out(o_16bit[8])
 );
 
m_not bi10 (
 .i_a(i_16bit[9]),
 .o_out(o_16bit[9])
 );
 
m_not bit11 (
 .i_a(i_16bit[10]),
 .o_out(o_16bit[10])
 );
 
m_not bit12 (
 .i_a(i_16bit[11]),
 .o_out(o_16bit[11])
 );
 
m_not bit13 (
 .i_a(i_16bit[12]),
 .o_out(o_16bit[12])
 );
 
m_not bit14 (
 .i_a(i_16bit[13]),
 .o_out(o_16bit[13])
 );
 
m_not bit15 (
 .i_a(i_16bit[14]),
 .o_out(o_16bit[14])
 );
 
m_not bit16 (
 .i_a(i_16bit[15]),
 .o_out(o_16bit[15])
 );
